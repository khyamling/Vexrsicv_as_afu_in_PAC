module bram_reset_in (
		input  wire  clk,         //       clk.clk
		input  wire  in_reset_n,  //  in_reset.reset_n
		output wire  out_reset_n  // out_reset.reset_n
	);
endmodule

